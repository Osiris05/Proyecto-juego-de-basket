��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  ����    Se�al (Clock)                    ���  CLED�� 	 CTerminal  ����        '����@��W8
IC=  �  ����        G����@��W8
IC�    ����        ��      �� 	 CResistor��  CValue  ����    180          �f@      �?   �  �p��               @P��O�HC=  �  ����        '����@P��O�HC�    ����         ��      �� 
 CPushBreak��  CKey  � J f         �  � d� y                 �|��H��  �  � 8� M                 �|��H�?    � L� d          ��    ��  �#�    10k          ��@      �?k  �  (x)�               @�, Օ3?  �  (�)�        =I.:V��?�, Օ3�    $�,�         ��      ��  CNPN��  CDummyValue  p�p�    100hFE            Y@      �? hFE �  p�q�         G����@���e>  �  H�]�        =I.:V��?�������  �  p�q�                 U�����    \�x�     #    ��      ��  K�k�    10k          ��@      �?k  �  phq}               @�e���>  �  p�q�        G����@�e����    l|t�     (    ��      ��  CBattery�  k �� �    3V(          @      �? V �  � �� �               @-�'h���  �  � �� 	                -�'h��?    � �� �     -    ��      �� 	 CIsolator�  ��         =I.:V��?��,Օ3?  �  � �� �         �<�e��?�|��H�?  �  � � !                �|��H��  �  !                 ��,Օ3�    � �     1  
 ��      ��  � �� �    100           Y@      �?   �  � x� �               @�|��H�?  �  � �� �        �<�e��?�|��H��    � �� �     7    ��                    ���  CWire  p���      :�  � �q�       :�  (`qa      :�  p`�a      :�  �`�q       :�  ����      :�  � �� �       :�  � x� �        :�  �  � 9       :�  8q9       :�  p8q�        :�  p�q9        :�   9        :�  (�)�       :�  (�)�       :�  (�I�      :�  �)�      :�  � `)a      :�  (`)y       :�  � `� y       :�  p`qi       :�  � `� a      :�  p�q�       :�  � � �        :�  � `� �       :�  � �� �                     �                              @  ;   ?    @   B  C   M    I # Q # $ J $ % % F ( O ( ) ) Q - S - . . R 1 K 1 2 T 2 3 3 C 4 4 G 7 N 7 8 8 T #  A E L O = ? >    R B  < 3  G F D < % E 4 D I K  J H $ 1 H N M =  P 7 > ( S L ) ; . A P - 8 2   +         �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 